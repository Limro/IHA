  --Example instantiation for system 'SOPC_System'
  SOPC_System_inst : SOPC_System
    port map(
      E_ci_multi_clock_from_the_cpu_0 => E_ci_multi_clock_from_the_cpu_0,
      E_ci_multi_reset_from_the_cpu_0 => E_ci_multi_reset_from_the_cpu_0,
      LCD_E_from_the_lcd_0 => LCD_E_from_the_lcd_0,
      LCD_RS_from_the_lcd_0 => LCD_RS_from_the_lcd_0,
      LCD_RW_from_the_lcd_0 => LCD_RW_from_the_lcd_0,
      LCD_data_to_and_from_the_lcd_0 => LCD_data_to_and_from_the_lcd_0,
      SRAM_ADDR_from_the_sram_0 => SRAM_ADDR_from_the_sram_0,
      SRAM_CE_N_from_the_sram_0 => SRAM_CE_N_from_the_sram_0,
      SRAM_DQ_to_and_from_the_sram_0 => SRAM_DQ_to_and_from_the_sram_0,
      SRAM_LB_N_from_the_sram_0 => SRAM_LB_N_from_the_sram_0,
      SRAM_OE_N_from_the_sram_0 => SRAM_OE_N_from_the_sram_0,
      SRAM_UB_N_from_the_sram_0 => SRAM_UB_N_from_the_sram_0,
      SRAM_WE_N_from_the_sram_0 => SRAM_WE_N_from_the_sram_0,
      clocks_0_sys_clk_out => clocks_0_sys_clk_out,
      hex0_from_the_mm_bus_seven_seg_four_digit_1 => hex0_from_the_mm_bus_seven_seg_four_digit_1,
      hex1_from_the_mm_bus_seven_seg_four_digit_1 => hex1_from_the_mm_bus_seven_seg_four_digit_1,
      hex2_from_the_mm_bus_seven_seg_four_digit_1 => hex2_from_the_mm_bus_seven_seg_four_digit_1,
      hex3_from_the_mm_bus_seven_seg_four_digit_1 => hex3_from_the_mm_bus_seven_seg_four_digit_1,
      out_port_from_the_pio_output_0 => out_port_from_the_pio_output_0,
      out_port_from_the_pio_output_1 => out_port_from_the_pio_output_1,
      clk_0 => clk_0,
      in_port_to_the_pio_input_0 => in_port_to_the_pio_input_0,
      reset_n => reset_n
    );


