  --Example instantiation for system 'CPU_System'
  CPU_System_inst : CPU_System
    port map(
      I2C_SCLK_from_the_audio_and_video_config_0 => I2C_SCLK_from_the_audio_and_video_config_0,
      I2C_SDAT_to_and_from_the_audio_and_video_config_0 => I2C_SDAT_to_and_from_the_audio_and_video_config_0,
      LCD_E_from_the_lcd_0 => LCD_E_from_the_lcd_0,
      LCD_RS_from_the_lcd_0 => LCD_RS_from_the_lcd_0,
      LCD_RW_from_the_lcd_0 => LCD_RW_from_the_lcd_0,
      LCD_data_to_and_from_the_lcd_0 => LCD_data_to_and_from_the_lcd_0,
      PS2_CLK_to_and_from_the_ps2_port => PS2_CLK_to_and_from_the_ps2_port,
      PS2_DAT_to_and_from_the_ps2_port => PS2_DAT_to_and_from_the_ps2_port,
      SRAM_ADDR_from_the_sram_0 => SRAM_ADDR_from_the_sram_0,
      SRAM_CE_N_from_the_sram_0 => SRAM_CE_N_from_the_sram_0,
      SRAM_DQ_to_and_from_the_sram_0 => SRAM_DQ_to_and_from_the_sram_0,
      SRAM_LB_N_from_the_sram_0 => SRAM_LB_N_from_the_sram_0,
      SRAM_OE_N_from_the_sram_0 => SRAM_OE_N_from_the_sram_0,
      SRAM_UB_N_from_the_sram_0 => SRAM_UB_N_from_the_sram_0,
      SRAM_WE_N_from_the_sram_0 => SRAM_WE_N_from_the_sram_0,
      dacdat_from_the_iis2st_0 => dacdat_from_the_iis2st_0,
      hex0_from_the_mm_bus_seven_seg_four_digit_0 => hex0_from_the_mm_bus_seven_seg_four_digit_0,
      hex1_from_the_mm_bus_seven_seg_four_digit_0 => hex1_from_the_mm_bus_seven_seg_four_digit_0,
      hex2_from_the_mm_bus_seven_seg_four_digit_0 => hex2_from_the_mm_bus_seven_seg_four_digit_0,
      hex3_from_the_mm_bus_seven_seg_four_digit_0 => hex3_from_the_mm_bus_seven_seg_four_digit_0,
      adcdat_to_the_iis2st_0 => adcdat_to_the_iis2st_0,
      adclrck_to_the_iis2st_0 => adclrck_to_the_iis2st_0,
      bitclk_to_the_iis2st_0 => bitclk_to_the_iis2st_0,
      clk_12 => clk_12,
      clk_50 => clk_50,
      daclrck_to_the_iis2st_0 => daclrck_to_the_iis2st_0,
      in_port_to_the_pio_input_key => in_port_to_the_pio_input_key,
      in_port_to_the_pio_input_sw => in_port_to_the_pio_input_sw,
      reset_n => reset_n
    );


