// mm_bus_seven_seg_four_digit_0.v

// Generated using ACDS version 12.1 177 at 2013.03.15.14:20:49

`timescale 1 ps / 1 ps
module mm_bus_seven_seg_four_digit_0 (
		input  wire        csi_clockreset_clk,     //       clockreset.clk
		input  wire        csi_clockreset_reset_n, // clockreset_reset.reset_n
		input  wire        avs_s1_write,           //               s1.write
		input  wire        avs_s1_read,            //                 .read
		input  wire        avs_s1_chipselect,      //                 .chipselect
		input  wire [7:0]  avs_s1_address,         //                 .address
		input  wire [15:0] avs_s1_writedata,       //                 .writedata
		output wire [15:0] avs_s1_readdata,        //                 .readdata
		output wire [6:0]  hex0,                   //              HEX.export
		output wire [6:0]  hex1,                   //                 .export
		output wire [6:0]  hex2,                   //                 .export
		output wire [6:0]  hex3                    //                 .export
	);

	mm_bus_seven_seg_four_digit mm_bus_seven_seg_four_digit_0_inst (
		.csi_clockreset_clk     (csi_clockreset_clk),     //       clockreset.clk
		.csi_clockreset_reset_n (csi_clockreset_reset_n), // clockreset_reset.reset_n
		.avs_s1_write           (avs_s1_write),           //               s1.write
		.avs_s1_read            (avs_s1_read),            //                 .read
		.avs_s1_chipselect      (avs_s1_chipselect),      //                 .chipselect
		.avs_s1_address         (avs_s1_address),         //                 .address
		.avs_s1_writedata       (avs_s1_writedata),       //                 .writedata
		.avs_s1_readdata        (avs_s1_readdata),        //                 .readdata
		.hex0                   (hex0),                   //              HEX.export
		.hex1                   (hex1),                   //                 .export
		.hex2                   (hex2),                   //                 .export
		.hex3                   (hex3)                    //                 .export
	);

endmodule
