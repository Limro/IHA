// FIRFilter_hw_0.v

// Generated using ACDS version 12.1 177 at 2013.03.06.11:37:31

`timescale 1 ps / 1 ps
module FIRFilter_hw_0 (
		input  wire        clk,              //                   clock.clk
		input  wire        reset_n,          //                   reset.reset_n
		input  wire [23:0] ast_sink_data,    //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,   //                        .valid
		input  wire [1:0]  ast_sink_error,   //                        .error
		input  wire        ast_sink_ready,   //                        .ready
		output wire [23:0] ast_source_data,  // avalon_streaming_source.data
		output wire        ast_source_valid, //                        .valid
		output wire [1:0]  ast_source_error, //                        .error
		output wire        ast_source_ready  //                        .ready
	);

	Fir firfilter_hw_0_inst (
		.clk              (clk),              //                   clock.clk
		.reset_n          (reset_n),          //                   reset.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_sink_ready   (ast_sink_ready),   //                        .ready
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error), //                        .error
		.ast_source_ready (ast_source_ready)  //                        .ready
	);

endmodule
